`uvm_analysis_imp_decl(_mon_cg)

class alu_coverage extends uvm_component;
  alu_sequence_item t1,t2;
  real drv1_cov,mon1_cov;
  `uvm_component_utils(alu_coverage)
  
  uvm_analysis_imp_mon_cg #(alu_sequence_item, alu_coverage) cov_mon;

  
  covergroup monitor_cov;
    ERR      : coverpoint t2.ERR {bins err[]={0,1};}
    COUT     : coverpoint t2.COUT {bins cout[]={0,1};}
    OFLOW    : coverpoint t2.OFLOW {bins oflow[]={0,1};}
    E        : coverpoint t2.E {bins e[]={0,1};}
    G        : coverpoint t2.G {bins g[]={0,1};}
    L        : coverpoint t2.L {bins l[]={0,1};}
    RES      : coverpoint t2.RES {bins res[]={[0:(1<<(`N+1))-1]};}
                                                
  endgroup
  
   function new(string name="alu_coverage",uvm_component parent);
    super.new(name,parent);
    cov_mon=new("cov_mon",this);
    cov_dri=new("cov_dri",this);
    driver_cov=new;
    monitor_cov=new;
  endfunction
    
   function void write_mon_cg(alu_sequence_item t);
    t2 = t;
    monitor_cov.sample();
     `uvm_info(get_type_name(),$sformatf("DATA RECEIVED FROM MONITOR IN COV,ERR=%d,OFLOW=%d,COUT=%d,E=%d,G=%d,L=%d,RES=%d",t2.ERR,t2.OFLOW,t2.COUT,t2.E,t2.G,t2.L,t2.RES),UVM_NONE);
  endfunction
  
   function void extract_phase(uvm_phase phase);
     super.extract_phase(phase);
    mon1_cov = monitor_cov.get_coverage();
  endfunction

  function void report_phase(uvm_phase phase);
    super.report_phase(phase);
    `uvm_info(get_type_name, $sformatf("[MONITOR] Coverage ------> %0.2f%%", mon1_cov), UVM_MEDIUM);
  endfunction
    
endclass
